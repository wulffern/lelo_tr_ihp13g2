magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741734000
<< checkpaint >>
rect 0 0 3168 1200
<< poly >>
rect 198 -40 330 40
rect 462 -40 594 40
rect 990 -40 1122 40
rect 1254 -40 1386 40
rect 1782 -40 1914 40
rect 2046 -40 2178 40
rect 2574 -40 2706 40
rect 2838 -40 2970 40
rect 198 40 330 120
rect 462 40 594 120
rect 990 40 1122 120
rect 1254 40 1386 120
rect 1782 40 1914 120
rect 2046 40 2178 120
rect 2574 40 2706 120
rect 2838 40 2970 120
rect 198 120 330 200
rect 462 120 594 200
rect 990 120 1122 200
rect 1254 120 1386 200
rect 1782 120 1914 200
rect 2046 120 2178 200
rect 2574 120 2706 200
rect 2838 120 2970 200
rect 198 840 330 920
rect 462 840 594 920
rect 990 840 1122 920
rect 1254 840 1386 920
rect 1782 840 1914 920
rect 2046 840 2178 920
rect 2574 840 2706 920
rect 2838 840 2970 920
rect 198 920 330 1000
rect 462 920 594 1000
rect 990 920 1122 1000
rect 1254 920 1386 1000
rect 1782 920 1914 1000
rect 2046 920 2178 1000
rect 2574 920 2706 1000
rect 2838 920 2970 1000
rect 198 1000 330 1080
rect 462 1000 594 1080
rect 990 1000 1122 1080
rect 1254 1000 1386 1080
rect 1782 1000 1914 1080
rect 2046 1000 2178 1080
rect 2574 1000 2706 1080
rect 2838 1000 2970 1080
rect -66 -40 66 40
rect 726 -40 858 40
rect 1518 -40 1650 40
rect 2310 -40 2442 40
rect 3102 -40 3234 40
rect -66 40 66 120
rect 726 40 858 120
rect 1518 40 1650 120
rect 2310 40 2442 120
rect 3102 40 3234 120
rect -66 120 66 200
rect 726 120 858 200
rect 1518 120 1650 200
rect 2310 120 2442 200
rect 3102 120 3234 200
rect -66 200 66 280
rect 726 200 858 280
rect 1518 200 1650 280
rect 2310 200 2442 280
rect 3102 200 3234 280
rect -66 280 66 360
rect 726 280 858 360
rect 1518 280 1650 360
rect 2310 280 2442 360
rect 3102 280 3234 360
rect -66 360 66 440
rect 726 360 858 440
rect 1518 360 1650 440
rect 2310 360 2442 440
rect 3102 360 3234 440
rect -66 440 66 520
rect 726 440 858 520
rect 1518 440 1650 520
rect 2310 440 2442 520
rect 3102 440 3234 520
rect -66 520 66 600
rect 726 520 858 600
rect 1518 520 1650 600
rect 2310 520 2442 600
rect 3102 520 3234 600
rect -66 600 66 680
rect 726 600 858 680
rect 1518 600 1650 680
rect 2310 600 2442 680
rect 3102 600 3234 680
rect -66 680 66 760
rect 726 680 858 760
rect 1518 680 1650 760
rect 2310 680 2442 760
rect 3102 680 3234 760
rect -66 760 66 840
rect 726 760 858 840
rect 1518 760 1650 840
rect 2310 760 2442 840
rect 3102 760 3234 840
rect -66 840 66 920
rect 726 840 858 920
rect 1518 840 1650 920
rect 2310 840 2442 920
rect 3102 840 3234 920
rect -66 920 66 1000
rect 726 920 858 1000
rect 1518 920 1650 1000
rect 2310 920 2442 1000
rect 3102 920 3234 1000
rect -66 1000 66 1080
rect 726 1000 858 1080
rect 1518 1000 1650 1080
rect 2310 1000 2442 1080
rect 3102 1000 3234 1080
<< xpolyres >>
rect 198 200 330 280
rect 462 200 594 280
rect 990 200 1122 280
rect 1254 200 1386 280
rect 1782 200 1914 280
rect 2046 200 2178 280
rect 2574 200 2706 280
rect 2838 200 2970 280
rect 198 280 330 360
rect 462 280 594 360
rect 990 280 1122 360
rect 1254 280 1386 360
rect 1782 280 1914 360
rect 2046 280 2178 360
rect 2574 280 2706 360
rect 2838 280 2970 360
rect 198 360 330 440
rect 462 360 594 440
rect 990 360 1122 440
rect 1254 360 1386 440
rect 1782 360 1914 440
rect 2046 360 2178 440
rect 2574 360 2706 440
rect 2838 360 2970 440
rect 198 440 330 520
rect 462 440 594 520
rect 990 440 1122 520
rect 1254 440 1386 520
rect 1782 440 1914 520
rect 2046 440 2178 520
rect 2574 440 2706 520
rect 2838 440 2970 520
rect 198 520 330 600
rect 462 520 594 600
rect 990 520 1122 600
rect 1254 520 1386 600
rect 1782 520 1914 600
rect 2046 520 2178 600
rect 2574 520 2706 600
rect 2838 520 2970 600
rect 198 600 330 680
rect 462 600 594 680
rect 990 600 1122 680
rect 1254 600 1386 680
rect 1782 600 1914 680
rect 2046 600 2178 680
rect 2574 600 2706 680
rect 2838 600 2970 680
rect 198 680 330 760
rect 462 680 594 760
rect 990 680 1122 760
rect 1254 680 1386 760
rect 1782 680 1914 760
rect 2046 680 2178 760
rect 2574 680 2706 760
rect 2838 680 2970 760
rect 198 760 330 840
rect 462 760 594 840
rect 990 760 1122 840
rect 1254 760 1386 840
rect 1782 760 1914 840
rect 2046 760 2178 840
rect 2574 760 2706 840
rect 2838 760 2970 840
<< pc >>
rect 231 40 297 80
rect 231 80 297 120
rect 495 40 561 80
rect 495 80 561 120
rect 1023 40 1089 80
rect 1023 80 1089 120
rect 1287 40 1353 80
rect 1287 80 1353 120
rect 1815 40 1881 80
rect 1815 80 1881 120
rect 2079 40 2145 80
rect 2079 80 2145 120
rect 2607 40 2673 80
rect 2607 80 2673 120
rect 2871 40 2937 80
rect 2871 80 2937 120
rect 231 920 297 960
rect 231 960 297 1000
rect 495 920 561 960
rect 495 960 561 1000
rect 1023 920 1089 960
rect 1023 960 1089 1000
rect 1287 920 1353 960
rect 1287 960 1353 1000
rect 1815 920 1881 960
rect 1815 960 1881 1000
rect 2079 920 2145 960
rect 2079 960 2145 1000
rect 2607 920 2673 960
rect 2607 960 2673 1000
rect 2871 920 2937 960
rect 2871 960 2937 1000
<< metal1 >>
rect 198 -40 594 40
rect 990 -40 1386 40
rect 1782 -40 2178 40
rect 2574 -40 2970 40
rect 198 40 594 120
rect 990 40 1386 120
rect 1782 40 2178 120
rect 2574 40 2970 120
rect 198 120 594 200
rect 990 120 1386 200
rect 1782 120 2178 200
rect 2574 120 2970 200
rect 198 840 330 920
rect 462 840 594 920
rect 990 840 1122 920
rect 1254 840 1386 920
rect 1782 840 1914 920
rect 2046 840 2178 920
rect 2574 840 2706 920
rect 2838 840 2970 920
rect 198 920 330 1000
rect 462 920 594 1000
rect 990 920 1122 1000
rect 1254 920 1386 1000
rect 1782 920 1914 1000
rect 2046 920 2178 1000
rect 2574 920 2706 1000
rect 2838 920 2970 1000
rect 198 1000 330 1080
rect 462 1000 594 1080
rect 990 1000 1122 1080
rect 1254 1000 1386 1080
rect 1782 1000 1914 1080
rect 2046 1000 2178 1080
rect 2574 1000 2706 1080
rect 2838 1000 2970 1080
rect 198 1080 330 1160
rect 462 1080 594 1160
rect 990 1080 1122 1160
rect 1254 1080 1386 1160
rect 1782 1080 1914 1160
rect 2046 1080 2178 1160
rect 2574 1080 2706 1160
rect 2838 1080 2970 1160
rect -66 1160 330 1240
rect -66 1160 330 1240
rect 462 1160 1122 1240
rect 2838 1160 3234 1240
rect 1254 1160 1914 1240
rect 2046 1160 2706 1240
rect 2838 1160 3234 1240
<< pwell >>
rect -66 -40 3234 1240
<< labels >>
flabel metal1 s -66 1160 330 1240 0 FreeSans 400 0 0 0 N
port 1 nsew signal bidirectional
flabel metal1 s 2838 1160 3234 1240 0 FreeSans 400 0 0 0 P
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 3168 1200
<< end >>
