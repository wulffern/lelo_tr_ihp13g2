magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741734000
<< checkpaint >>
rect 0 0 3728 1760
<< metal1 >>
rect 16 16 3712 128
rect 128 16 3600 128
rect 16 16 3712 128
rect 128 1632 3600 1744
rect 16 1632 3712 1744
rect 16 128 128 1632
rect 16 16 128 1744
rect 3600 128 3712 1632
rect 3600 16 3712 1744
rect 16 16 3712 128
rect 3118 1440 3514 1520
rect 214 1440 610 1520
<< ptapc >>
rect 144 32 224 112
rect 224 32 304 112
rect 304 32 384 112
rect 384 32 464 112
rect 464 32 544 112
rect 544 32 624 112
rect 624 32 704 112
rect 704 32 784 112
rect 784 32 864 112
rect 864 32 944 112
rect 944 32 1024 112
rect 1024 32 1104 112
rect 1104 32 1184 112
rect 1184 32 1264 112
rect 1264 32 1344 112
rect 1344 32 1424 112
rect 1424 32 1504 112
rect 1504 32 1584 112
rect 1584 32 1664 112
rect 1664 32 1744 112
rect 1744 32 1824 112
rect 1824 32 1904 112
rect 1904 32 1984 112
rect 1984 32 2064 112
rect 2064 32 2144 112
rect 2144 32 2224 112
rect 2224 32 2304 112
rect 2304 32 2384 112
rect 2384 32 2464 112
rect 2464 32 2544 112
rect 2544 32 2624 112
rect 2624 32 2704 112
rect 2704 32 2784 112
rect 2784 32 2864 112
rect 2864 32 2944 112
rect 2944 32 3024 112
rect 3024 32 3104 112
rect 3104 32 3184 112
rect 3184 32 3264 112
rect 3264 32 3344 112
rect 3344 32 3424 112
rect 3424 32 3504 112
rect 3504 32 3584 112
rect 144 1648 224 1728
rect 224 1648 304 1728
rect 304 1648 384 1728
rect 384 1648 464 1728
rect 464 1648 544 1728
rect 544 1648 624 1728
rect 624 1648 704 1728
rect 704 1648 784 1728
rect 784 1648 864 1728
rect 864 1648 944 1728
rect 944 1648 1024 1728
rect 1024 1648 1104 1728
rect 1104 1648 1184 1728
rect 1184 1648 1264 1728
rect 1264 1648 1344 1728
rect 1344 1648 1424 1728
rect 1424 1648 1504 1728
rect 1504 1648 1584 1728
rect 1584 1648 1664 1728
rect 1664 1648 1744 1728
rect 1744 1648 1824 1728
rect 1824 1648 1904 1728
rect 1904 1648 1984 1728
rect 1984 1648 2064 1728
rect 2064 1648 2144 1728
rect 2144 1648 2224 1728
rect 2224 1648 2304 1728
rect 2304 1648 2384 1728
rect 2384 1648 2464 1728
rect 2464 1648 2544 1728
rect 2544 1648 2624 1728
rect 2624 1648 2704 1728
rect 2704 1648 2784 1728
rect 2784 1648 2864 1728
rect 2864 1648 2944 1728
rect 2944 1648 3024 1728
rect 3024 1648 3104 1728
rect 3104 1648 3184 1728
rect 3184 1648 3264 1728
rect 3264 1648 3344 1728
rect 3344 1648 3424 1728
rect 3424 1648 3504 1728
rect 3504 1648 3584 1728
rect 32 160 112 240
rect 32 240 112 320
rect 32 320 112 400
rect 32 400 112 480
rect 32 480 112 560
rect 32 560 112 640
rect 32 640 112 720
rect 32 720 112 800
rect 32 800 112 880
rect 32 880 112 960
rect 32 960 112 1040
rect 32 1040 112 1120
rect 32 1120 112 1200
rect 32 1200 112 1280
rect 32 1280 112 1360
rect 32 1360 112 1440
rect 32 1440 112 1520
rect 32 1520 112 1600
rect 3616 160 3696 240
rect 3616 240 3696 320
rect 3616 320 3696 400
rect 3616 400 3696 480
rect 3616 480 3696 560
rect 3616 560 3696 640
rect 3616 640 3696 720
rect 3616 720 3696 800
rect 3616 800 3696 880
rect 3616 880 3696 960
rect 3616 960 3696 1040
rect 3616 1040 3696 1120
rect 3616 1120 3696 1200
rect 3616 1200 3696 1280
rect 3616 1280 3696 1360
rect 3616 1360 3696 1440
rect 3616 1440 3696 1520
rect 3616 1520 3696 1600
<< ptap >>
rect 0 0 3728 144
rect 0 1616 3728 1760
rect 0 0 144 1760
rect 3584 0 3728 1760
use LELOTR_RES8 XA1 
transform 1 0 280 0 1 280
box 280 280 3448 1480
<< labels >>
flabel metal1 s 16 16 3712 128 0 FreeSans 400 0 0 0 B
port 3 nsew signal bidirectional
flabel metal1 s 3118 1440 3514 1520 0 FreeSans 400 0 0 0 P
port 1 nsew signal bidirectional
flabel metal1 s 214 1440 610 1520 0 FreeSans 400 0 0 0 N
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 3728 1760
<< end >>
