magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741734000
<< checkpaint >>
rect 0 0 1628 320
<< metal1 >>
rect -66 140 374 180
rect 286 140 418 180
rect 418 60 594 100
rect 418 60 458 180
rect 286 140 418 180
rect 418 220 594 260
rect 418 140 458 260
rect 1034 60 1166 100
rect 1166 140 1342 180
rect 1166 60 1206 180
rect 1034 220 1166 260
rect 1166 140 1342 180
rect 1166 140 1206 260
rect 1254 140 1694 180
<< metal4 >>
rect 946 0 1098 320
rect 506 0 658 320
rect 946 0 1098 320
rect 506 0 658 320
use LELOTR_NCHDL MN1 
transform 1 0 0 0 1 0
box 0 0 814 320
use LELOTR_PCHDL MP1 
transform 1 0 814 0 1 0
box 814 0 1628 320
use LELOTR_cut_M1M4_2x1 xcut0 
transform 1 0 946 0 1 220
box 946 220 1098 262
use LELOTR_cut_M1M4_2x1 xcut1 
transform 1 0 946 0 1 60
box 946 60 1098 102
use LELOTR_cut_M1M4_2x1 xcut2 
transform 1 0 506 0 1 220
box 506 220 658 262
use LELOTR_cut_M1M4_2x1 xcut3 
transform 1 0 506 0 1 60
box 506 60 658 102
<< labels >>
flabel metal4 s 946 0 1098 320 0 FreeSans 400 0 0 0 AVDD
port 1 nsew signal bidirectional
flabel metal4 s 506 0 658 320 0 FreeSans 400 0 0 0 AVSS
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1628 320
<< end >>
