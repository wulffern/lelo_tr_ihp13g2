magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741734000
<< checkpaint >>
rect 0 0 1628 480
<< metal1 >>
rect 594 380 726 420
rect 726 220 1034 260
rect 726 220 766 420
rect 574 220 614 260
rect 198 140 374 180
rect 198 300 374 340
rect 506 380 682 420
<< poly >>
rect 242 146 1386 174
rect 242 306 1386 334
<< metal4 >>
rect 946 0 1098 480
rect 506 0 658 480
rect 946 0 1098 480
rect 506 0 658 480
use LELOTR_NCHDL MN0 
transform 1 0 0 0 1 0
box 0 0 814 320
use LELOTR_NCHDL MN1 
transform 1 0 0 0 1 160
box 0 160 814 480
use LELOTR_PCHDL MP0 
transform 1 0 814 0 1 0
box 814 0 1628 320
use LELOTR_PCHDL MP1 
transform 1 0 814 0 1 160
box 814 160 1628 480
use LELOTR_cut_M1M4_2x1 xcut0 
transform 1 0 946 0 1 60
box 946 60 1098 102
use LELOTR_cut_M1M4_2x1 xcut1 
transform 1 0 946 0 1 380
box 946 380 1098 422
use LELOTR_cut_M1M4_2x1 xcut2 
transform 1 0 506 0 1 60
box 506 60 658 102
<< labels >>
flabel metal1 s 198 140 374 180 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel metal1 s 198 300 374 340 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
flabel metal1 s 506 380 682 420 0 FreeSans 400 0 0 0 Y
port 3 nsew signal bidirectional
flabel metal4 s 946 0 1098 480 0 FreeSans 400 0 0 0 AVDD
port 4 nsew signal bidirectional
flabel metal4 s 506 0 658 480 0 FreeSans 400 0 0 0 AVSS
port 5 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1628 480
<< end >>
