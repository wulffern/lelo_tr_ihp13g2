magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741993200
<< checkpaint >>
rect 0 0 1628 640
<< metal1 >>
rect 594 60 726 100
rect 726 60 1034 100
rect 726 60 766 100
rect 594 540 726 580
rect 726 540 1034 580
rect 726 540 766 580
rect 594 380 726 420
rect 726 380 1034 420
rect 726 380 766 420
rect 266 140 306 340
rect 286 460 418 500
rect 418 60 594 100
rect 418 60 458 500
rect 1342 140 1474 180
rect 1342 460 1474 500
rect 1474 140 1514 500
rect 1034 220 1166 260
rect 1166 300 1342 340
rect 1166 220 1206 340
rect 1254 140 1430 180
rect 946 380 1122 420
rect 506 540 682 580
<< poly >>
rect 242 146 1386 174
<< metal4 >>
rect 946 0 1098 640
rect 506 0 658 640
rect 946 0 1098 640
rect 506 0 658 640
use LELOTR_NCHDL MN0 
transform 1 0 0 0 1 0
box 0 0 814 320
use LELOTR_NCHDL MN1 
transform 1 0 0 0 1 160
box 0 160 814 480
use LELOTR_NCHDL MN2 
transform 1 0 0 0 1 320
box 0 320 814 640
use LELOTR_PCHDL MP0 
transform 1 0 814 0 1 0
box 814 0 1628 320
use LELOTR_PCHDL MP1_DMY 
transform 1 0 814 0 1 160
box 814 160 1628 480
use LELOTR_PCHDL MP2 
transform 1 0 814 0 1 320
box 814 320 1628 640
use LELOTR_cut_M1M4_2x1 xcut0 
transform 1 0 946 0 1 220
box 946 220 1098 262
use LELOTR_cut_M1M4_2x1 xcut1 
transform 1 0 506 0 1 220
box 506 220 658 262
use LELOTR_cut_M1M4_2x1 xcut2 
transform 1 0 506 0 1 220
box 506 220 658 262
<< labels >>
flabel metal1 s 1254 140 1430 180 0 FreeSans 400 0 0 0 C
port 1 nsew signal bidirectional
flabel metal1 s 946 380 1122 420 0 FreeSans 400 0 0 0 B
port 3 nsew signal bidirectional
flabel metal1 s 506 540 682 580 0 FreeSans 400 0 0 0 A
port 2 nsew signal bidirectional
flabel metal4 s 946 0 1098 640 0 FreeSans 400 0 0 0 AVDD
port 4 nsew signal bidirectional
flabel metal4 s 506 0 658 640 0 FreeSans 400 0 0 0 AVSS
port 5 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1628 640
<< end >>
