
*.subckt CAPX1 A B
*C1 B A sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
*.ends
