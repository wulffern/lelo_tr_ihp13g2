magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741734000
<< checkpaint >>
rect 0 0 1352 1760
<< metal1 >>
rect 16 16 1336 128
rect 128 16 1224 128
rect 16 16 1336 128
rect 128 1632 1224 1744
rect 16 1632 1336 1744
rect 16 128 128 1632
rect 16 16 128 1744
rect 1224 128 1336 1632
rect 1224 16 1336 1744
rect 16 16 1336 128
rect 742 1440 1138 1520
rect 214 1440 610 1520
<< ptapc >>
rect 156 32 236 112
rect 236 32 316 112
rect 316 32 396 112
rect 396 32 476 112
rect 476 32 556 112
rect 556 32 636 112
rect 636 32 716 112
rect 716 32 796 112
rect 796 32 876 112
rect 876 32 956 112
rect 956 32 1036 112
rect 1036 32 1116 112
rect 1116 32 1196 112
rect 156 1648 236 1728
rect 236 1648 316 1728
rect 316 1648 396 1728
rect 396 1648 476 1728
rect 476 1648 556 1728
rect 556 1648 636 1728
rect 636 1648 716 1728
rect 716 1648 796 1728
rect 796 1648 876 1728
rect 876 1648 956 1728
rect 956 1648 1036 1728
rect 1036 1648 1116 1728
rect 1116 1648 1196 1728
rect 32 160 112 240
rect 32 240 112 320
rect 32 320 112 400
rect 32 400 112 480
rect 32 480 112 560
rect 32 560 112 640
rect 32 640 112 720
rect 32 720 112 800
rect 32 800 112 880
rect 32 880 112 960
rect 32 960 112 1040
rect 32 1040 112 1120
rect 32 1120 112 1200
rect 32 1200 112 1280
rect 32 1280 112 1360
rect 32 1360 112 1440
rect 32 1440 112 1520
rect 32 1520 112 1600
rect 1240 160 1320 240
rect 1240 240 1320 320
rect 1240 320 1320 400
rect 1240 400 1320 480
rect 1240 480 1320 560
rect 1240 560 1320 640
rect 1240 640 1320 720
rect 1240 720 1320 800
rect 1240 800 1320 880
rect 1240 880 1320 960
rect 1240 960 1320 1040
rect 1240 1040 1320 1120
rect 1240 1120 1320 1200
rect 1240 1200 1320 1280
rect 1240 1280 1320 1360
rect 1240 1360 1320 1440
rect 1240 1440 1320 1520
rect 1240 1520 1320 1600
<< ptap >>
rect 0 0 1352 144
rect 0 1616 1352 1760
rect 0 0 144 1760
rect 1208 0 1352 1760
use LELOTR_RES2 XA1 
transform 1 0 280 0 1 280
box 280 280 1072 1480
<< labels >>
flabel metal1 s 16 16 1336 128 0 FreeSans 400 0 0 0 B
port 3 nsew signal bidirectional
flabel metal1 s 742 1440 1138 1520 0 FreeSans 400 0 0 0 P
port 1 nsew signal bidirectional
flabel metal1 s 214 1440 610 1520 0 FreeSans 400 0 0 0 N
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1352 1760
<< end >>
