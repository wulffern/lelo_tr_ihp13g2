magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741734000
<< checkpaint >>
rect 0 0 1628 1600
<< metal1 >>
rect 594 220 726 260
rect 594 380 726 420
rect 594 700 726 740
rect 594 1020 726 1060
rect 726 220 766 1060
rect 862 220 1034 260
rect 862 380 1034 420
rect 862 860 1034 900
rect 862 1180 1034 1220
rect 862 220 902 1220
rect 266 140 306 500
rect 1342 780 1474 820
rect 1082 580 1474 620
rect 1390 1140 1474 1180
rect 1390 1460 1474 1500
rect 1474 580 1514 1500
rect 1034 540 1122 580
rect 1342 1100 1430 1140
rect 1342 1420 1430 1460
rect 114 780 286 820
rect 114 580 546 620
rect 114 1140 238 1180
rect 114 1460 238 1500
rect 114 580 154 1500
rect 506 540 594 580
rect 198 1100 286 1140
rect 198 1420 286 1460
rect 422 860 594 900
rect 422 1180 594 1220
rect 422 860 462 1220
rect 594 1500 726 1540
rect 726 1500 1034 1540
rect 726 1500 766 1540
rect 594 1180 726 1220
rect 726 1340 1034 1380
rect 726 1180 766 1380
rect 1034 700 1166 740
rect 1034 1020 1166 1060
rect 1166 700 1206 1060
rect 198 140 374 180
rect 506 1500 682 1540
<< metal2 >>
rect 594 1340 726 1380
rect 726 1020 1034 1060
rect 726 1020 766 1380
rect 594 540 726 580
rect 726 540 1034 580
rect 726 540 766 580
<< poly >>
rect 242 146 1386 174
rect 242 466 1386 494
<< metal4 >>
rect 946 0 1098 1600
rect 506 0 658 1600
rect 946 0 1098 1600
rect 506 0 658 1600
use LELOTR_NCHDL XA2 
transform 1 0 0 0 1 0
box 0 0 814 320
use LELOTR_NCHDL XA3 
transform 1 0 0 0 1 320
box 0 320 814 640
use LELOTR_NCHDL XA4a 
transform 1 0 0 0 1 640
box 0 640 814 960
use LELOTR_NCHDL XA4b 
transform 1 0 0 0 1 960
box 0 960 814 1280
use LELOTR_NCHDL XA5 
transform 1 0 0 0 1 1280
box 0 1280 814 1600
use LELOTR_PCHDL XB0 
transform 1 0 814 0 1 0
box 814 0 1628 320
use LELOTR_PCHDL XB1 
transform 1 0 814 0 1 320
box 814 320 1628 640
use LELOTR_PCHDL XB3a 
transform 1 0 814 0 1 640
box 814 640 1628 960
use LELOTR_PCHDL XB3b 
transform 1 0 814 0 1 960
box 814 960 1628 1280
use LELOTR_PCHDL XB4 
transform 1 0 814 0 1 1280
box 814 1280 1628 1600
use LELOTR_cut_M1M2_2x1 xcut0 
transform 1 0 506 0 1 1340
box 506 1340 658 1382
use LELOTR_cut_M1M2_2x1 xcut1 
transform 1 0 946 0 1 1020
box 946 1020 1098 1062
use LELOTR_cut_M1M2_2x1 xcut2 
transform 1 0 506 0 1 540
box 506 540 658 582
use LELOTR_cut_M1M2_2x1 xcut3 
transform 1 0 946 0 1 540
box 946 540 1098 582
use LELOTR_cut_M1M4_2x1 xcut4 
transform 1 0 946 0 1 60
box 946 60 1098 102
use LELOTR_cut_M1M4_2x1 xcut5 
transform 1 0 946 0 1 1340
box 946 1340 1098 1382
use LELOTR_cut_M1M4_2x1 xcut6 
transform 1 0 506 0 1 60
box 506 60 658 102
use LELOTR_cut_M1M4_2x1 xcut7 
transform 1 0 506 0 1 1340
box 506 1340 658 1382
<< labels >>
flabel metal1 s 198 140 374 180 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel metal1 s 506 1500 682 1540 0 FreeSans 400 0 0 0 Y
port 2 nsew signal bidirectional
flabel metal4 s 946 0 1098 1600 0 FreeSans 400 0 0 0 AVDD
port 3 nsew signal bidirectional
flabel metal4 s 506 0 658 1600 0 FreeSans 400 0 0 0 AVSS
port 4 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1628 1600
<< end >>
