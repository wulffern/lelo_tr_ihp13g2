magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741993200
<< checkpaint >>
rect 0 0 1584 1200
<< poly >>
rect 198 -40 330 40
rect 462 -40 594 40
rect 990 -40 1122 40
rect 1254 -40 1386 40
rect 198 40 330 120
rect 462 40 594 120
rect 990 40 1122 120
rect 1254 40 1386 120
rect 198 120 330 200
rect 462 120 594 200
rect 990 120 1122 200
rect 1254 120 1386 200
rect 198 840 330 920
rect 462 840 594 920
rect 990 840 1122 920
rect 1254 840 1386 920
rect 198 920 330 1000
rect 462 920 594 1000
rect 990 920 1122 1000
rect 1254 920 1386 1000
rect 198 1000 330 1080
rect 462 1000 594 1080
rect 990 1000 1122 1080
rect 1254 1000 1386 1080
rect -66 -40 66 40
rect 726 -40 858 40
rect 1518 -40 1650 40
rect -66 40 66 120
rect 726 40 858 120
rect 1518 40 1650 120
rect -66 120 66 200
rect 726 120 858 200
rect 1518 120 1650 200
rect -66 200 66 280
rect 726 200 858 280
rect 1518 200 1650 280
rect -66 280 66 360
rect 726 280 858 360
rect 1518 280 1650 360
rect -66 360 66 440
rect 726 360 858 440
rect 1518 360 1650 440
rect -66 440 66 520
rect 726 440 858 520
rect 1518 440 1650 520
rect -66 520 66 600
rect 726 520 858 600
rect 1518 520 1650 600
rect -66 600 66 680
rect 726 600 858 680
rect 1518 600 1650 680
rect -66 680 66 760
rect 726 680 858 760
rect 1518 680 1650 760
rect -66 760 66 840
rect 726 760 858 840
rect 1518 760 1650 840
rect -66 840 66 920
rect 726 840 858 920
rect 1518 840 1650 920
rect -66 920 66 1000
rect 726 920 858 1000
rect 1518 920 1650 1000
rect -66 1000 66 1080
rect 726 1000 858 1080
rect 1518 1000 1650 1080
<< xpolyres >>
rect 198 200 330 280
rect 462 200 594 280
rect 990 200 1122 280
rect 1254 200 1386 280
rect 198 280 330 360
rect 462 280 594 360
rect 990 280 1122 360
rect 1254 280 1386 360
rect 198 360 330 440
rect 462 360 594 440
rect 990 360 1122 440
rect 1254 360 1386 440
rect 198 440 330 520
rect 462 440 594 520
rect 990 440 1122 520
rect 1254 440 1386 520
rect 198 520 330 600
rect 462 520 594 600
rect 990 520 1122 600
rect 1254 520 1386 600
rect 198 600 330 680
rect 462 600 594 680
rect 990 600 1122 680
rect 1254 600 1386 680
rect 198 680 330 760
rect 462 680 594 760
rect 990 680 1122 760
rect 1254 680 1386 760
rect 198 760 330 840
rect 462 760 594 840
rect 990 760 1122 840
rect 1254 760 1386 840
<< pc >>
rect 231 40 297 80
rect 231 80 297 120
rect 495 40 561 80
rect 495 80 561 120
rect 1023 40 1089 80
rect 1023 80 1089 120
rect 1287 40 1353 80
rect 1287 80 1353 120
rect 231 920 297 960
rect 231 960 297 1000
rect 495 920 561 960
rect 495 960 561 1000
rect 1023 920 1089 960
rect 1023 960 1089 1000
rect 1287 920 1353 960
rect 1287 960 1353 1000
<< metal1 >>
rect 198 -40 594 40
rect 990 -40 1386 40
rect 198 40 594 120
rect 990 40 1386 120
rect 198 120 594 200
rect 990 120 1386 200
rect 198 840 330 920
rect 462 840 594 920
rect 990 840 1122 920
rect 1254 840 1386 920
rect 198 920 330 1000
rect 462 920 594 1000
rect 990 920 1122 1000
rect 1254 920 1386 1000
rect 198 1000 330 1080
rect 462 1000 594 1080
rect 990 1000 1122 1080
rect 1254 1000 1386 1080
rect 198 1080 330 1160
rect 462 1080 594 1160
rect 990 1080 1122 1160
rect 1254 1080 1386 1160
rect -66 1160 330 1240
rect -66 1160 330 1240
rect 462 1160 1122 1240
rect 1254 1160 1650 1240
rect 1254 1160 1650 1240
<< pwell >>
rect -66 -40 1650 1240
<< labels >>
flabel metal1 s -66 1160 330 1240 0 FreeSans 400 0 0 0 N
port 1 nsew signal bidirectional
flabel metal1 s 1254 1160 1650 1240 0 FreeSans 400 0 0 0 P
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1584 1200
<< end >>
