magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741734000
<< checkpaint >>
rect 0 0 6896 1760
<< metal1 >>
rect 16 16 6880 128
rect 128 16 6768 128
rect 16 16 6880 128
rect 128 1632 6768 1744
rect 16 1632 6880 1744
rect 16 128 128 1632
rect 16 16 128 1744
rect 6768 128 6880 1632
rect 6768 16 6880 1744
rect 16 16 6880 128
rect 6286 1440 6682 1520
rect 214 1440 610 1520
<< ptapc >>
rect 168 32 248 112
rect 248 32 328 112
rect 328 32 408 112
rect 408 32 488 112
rect 488 32 568 112
rect 568 32 648 112
rect 648 32 728 112
rect 728 32 808 112
rect 808 32 888 112
rect 888 32 968 112
rect 968 32 1048 112
rect 1048 32 1128 112
rect 1128 32 1208 112
rect 1208 32 1288 112
rect 1288 32 1368 112
rect 1368 32 1448 112
rect 1448 32 1528 112
rect 1528 32 1608 112
rect 1608 32 1688 112
rect 1688 32 1768 112
rect 1768 32 1848 112
rect 1848 32 1928 112
rect 1928 32 2008 112
rect 2008 32 2088 112
rect 2088 32 2168 112
rect 2168 32 2248 112
rect 2248 32 2328 112
rect 2328 32 2408 112
rect 2408 32 2488 112
rect 2488 32 2568 112
rect 2568 32 2648 112
rect 2648 32 2728 112
rect 2728 32 2808 112
rect 2808 32 2888 112
rect 2888 32 2968 112
rect 2968 32 3048 112
rect 3048 32 3128 112
rect 3128 32 3208 112
rect 3208 32 3288 112
rect 3288 32 3368 112
rect 3368 32 3448 112
rect 3448 32 3528 112
rect 3528 32 3608 112
rect 3608 32 3688 112
rect 3688 32 3768 112
rect 3768 32 3848 112
rect 3848 32 3928 112
rect 3928 32 4008 112
rect 4008 32 4088 112
rect 4088 32 4168 112
rect 4168 32 4248 112
rect 4248 32 4328 112
rect 4328 32 4408 112
rect 4408 32 4488 112
rect 4488 32 4568 112
rect 4568 32 4648 112
rect 4648 32 4728 112
rect 4728 32 4808 112
rect 4808 32 4888 112
rect 4888 32 4968 112
rect 4968 32 5048 112
rect 5048 32 5128 112
rect 5128 32 5208 112
rect 5208 32 5288 112
rect 5288 32 5368 112
rect 5368 32 5448 112
rect 5448 32 5528 112
rect 5528 32 5608 112
rect 5608 32 5688 112
rect 5688 32 5768 112
rect 5768 32 5848 112
rect 5848 32 5928 112
rect 5928 32 6008 112
rect 6008 32 6088 112
rect 6088 32 6168 112
rect 6168 32 6248 112
rect 6248 32 6328 112
rect 6328 32 6408 112
rect 6408 32 6488 112
rect 6488 32 6568 112
rect 6568 32 6648 112
rect 6648 32 6728 112
rect 168 1648 248 1728
rect 248 1648 328 1728
rect 328 1648 408 1728
rect 408 1648 488 1728
rect 488 1648 568 1728
rect 568 1648 648 1728
rect 648 1648 728 1728
rect 728 1648 808 1728
rect 808 1648 888 1728
rect 888 1648 968 1728
rect 968 1648 1048 1728
rect 1048 1648 1128 1728
rect 1128 1648 1208 1728
rect 1208 1648 1288 1728
rect 1288 1648 1368 1728
rect 1368 1648 1448 1728
rect 1448 1648 1528 1728
rect 1528 1648 1608 1728
rect 1608 1648 1688 1728
rect 1688 1648 1768 1728
rect 1768 1648 1848 1728
rect 1848 1648 1928 1728
rect 1928 1648 2008 1728
rect 2008 1648 2088 1728
rect 2088 1648 2168 1728
rect 2168 1648 2248 1728
rect 2248 1648 2328 1728
rect 2328 1648 2408 1728
rect 2408 1648 2488 1728
rect 2488 1648 2568 1728
rect 2568 1648 2648 1728
rect 2648 1648 2728 1728
rect 2728 1648 2808 1728
rect 2808 1648 2888 1728
rect 2888 1648 2968 1728
rect 2968 1648 3048 1728
rect 3048 1648 3128 1728
rect 3128 1648 3208 1728
rect 3208 1648 3288 1728
rect 3288 1648 3368 1728
rect 3368 1648 3448 1728
rect 3448 1648 3528 1728
rect 3528 1648 3608 1728
rect 3608 1648 3688 1728
rect 3688 1648 3768 1728
rect 3768 1648 3848 1728
rect 3848 1648 3928 1728
rect 3928 1648 4008 1728
rect 4008 1648 4088 1728
rect 4088 1648 4168 1728
rect 4168 1648 4248 1728
rect 4248 1648 4328 1728
rect 4328 1648 4408 1728
rect 4408 1648 4488 1728
rect 4488 1648 4568 1728
rect 4568 1648 4648 1728
rect 4648 1648 4728 1728
rect 4728 1648 4808 1728
rect 4808 1648 4888 1728
rect 4888 1648 4968 1728
rect 4968 1648 5048 1728
rect 5048 1648 5128 1728
rect 5128 1648 5208 1728
rect 5208 1648 5288 1728
rect 5288 1648 5368 1728
rect 5368 1648 5448 1728
rect 5448 1648 5528 1728
rect 5528 1648 5608 1728
rect 5608 1648 5688 1728
rect 5688 1648 5768 1728
rect 5768 1648 5848 1728
rect 5848 1648 5928 1728
rect 5928 1648 6008 1728
rect 6008 1648 6088 1728
rect 6088 1648 6168 1728
rect 6168 1648 6248 1728
rect 6248 1648 6328 1728
rect 6328 1648 6408 1728
rect 6408 1648 6488 1728
rect 6488 1648 6568 1728
rect 6568 1648 6648 1728
rect 6648 1648 6728 1728
rect 32 160 112 240
rect 32 240 112 320
rect 32 320 112 400
rect 32 400 112 480
rect 32 480 112 560
rect 32 560 112 640
rect 32 640 112 720
rect 32 720 112 800
rect 32 800 112 880
rect 32 880 112 960
rect 32 960 112 1040
rect 32 1040 112 1120
rect 32 1120 112 1200
rect 32 1200 112 1280
rect 32 1280 112 1360
rect 32 1360 112 1440
rect 32 1440 112 1520
rect 32 1520 112 1600
rect 6784 160 6864 240
rect 6784 240 6864 320
rect 6784 320 6864 400
rect 6784 400 6864 480
rect 6784 480 6864 560
rect 6784 560 6864 640
rect 6784 640 6864 720
rect 6784 720 6864 800
rect 6784 800 6864 880
rect 6784 880 6864 960
rect 6784 960 6864 1040
rect 6784 1040 6864 1120
rect 6784 1120 6864 1200
rect 6784 1200 6864 1280
rect 6784 1280 6864 1360
rect 6784 1360 6864 1440
rect 6784 1440 6864 1520
rect 6784 1520 6864 1600
<< ptap >>
rect 0 0 6896 144
rect 0 1616 6896 1760
rect 0 0 144 1760
rect 6752 0 6896 1760
use LELOTR_RES16 XA1 
transform 1 0 280 0 1 280
box 280 280 6616 1480
<< labels >>
flabel metal1 s 16 16 6880 128 0 FreeSans 400 0 0 0 B
port 3 nsew signal bidirectional
flabel metal1 s 6286 1440 6682 1520 0 FreeSans 400 0 0 0 P
port 1 nsew signal bidirectional
flabel metal1 s 214 1440 610 1520 0 FreeSans 400 0 0 0 N
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 6896 1760
<< end >>
