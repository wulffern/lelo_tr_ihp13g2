magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741734000
<< checkpaint >>
rect 0 0 2144 1760
<< metal1 >>
rect 16 16 2128 128
rect 128 16 2016 128
rect 16 16 2128 128
rect 128 1632 2016 1744
rect 16 1632 2128 1744
rect 16 128 128 1632
rect 16 16 128 1744
rect 2016 128 2128 1632
rect 2016 16 2128 1744
rect 16 16 2128 128
rect 1534 1440 1930 1520
rect 214 1440 610 1520
<< ptapc >>
rect 152 32 232 112
rect 232 32 312 112
rect 312 32 392 112
rect 392 32 472 112
rect 472 32 552 112
rect 552 32 632 112
rect 632 32 712 112
rect 712 32 792 112
rect 792 32 872 112
rect 872 32 952 112
rect 952 32 1032 112
rect 1032 32 1112 112
rect 1112 32 1192 112
rect 1192 32 1272 112
rect 1272 32 1352 112
rect 1352 32 1432 112
rect 1432 32 1512 112
rect 1512 32 1592 112
rect 1592 32 1672 112
rect 1672 32 1752 112
rect 1752 32 1832 112
rect 1832 32 1912 112
rect 1912 32 1992 112
rect 152 1648 232 1728
rect 232 1648 312 1728
rect 312 1648 392 1728
rect 392 1648 472 1728
rect 472 1648 552 1728
rect 552 1648 632 1728
rect 632 1648 712 1728
rect 712 1648 792 1728
rect 792 1648 872 1728
rect 872 1648 952 1728
rect 952 1648 1032 1728
rect 1032 1648 1112 1728
rect 1112 1648 1192 1728
rect 1192 1648 1272 1728
rect 1272 1648 1352 1728
rect 1352 1648 1432 1728
rect 1432 1648 1512 1728
rect 1512 1648 1592 1728
rect 1592 1648 1672 1728
rect 1672 1648 1752 1728
rect 1752 1648 1832 1728
rect 1832 1648 1912 1728
rect 1912 1648 1992 1728
rect 32 160 112 240
rect 32 240 112 320
rect 32 320 112 400
rect 32 400 112 480
rect 32 480 112 560
rect 32 560 112 640
rect 32 640 112 720
rect 32 720 112 800
rect 32 800 112 880
rect 32 880 112 960
rect 32 960 112 1040
rect 32 1040 112 1120
rect 32 1120 112 1200
rect 32 1200 112 1280
rect 32 1280 112 1360
rect 32 1360 112 1440
rect 32 1440 112 1520
rect 32 1520 112 1600
rect 2032 160 2112 240
rect 2032 240 2112 320
rect 2032 320 2112 400
rect 2032 400 2112 480
rect 2032 480 2112 560
rect 2032 560 2112 640
rect 2032 640 2112 720
rect 2032 720 2112 800
rect 2032 800 2112 880
rect 2032 880 2112 960
rect 2032 960 2112 1040
rect 2032 1040 2112 1120
rect 2032 1120 2112 1200
rect 2032 1200 2112 1280
rect 2032 1280 2112 1360
rect 2032 1360 2112 1440
rect 2032 1440 2112 1520
rect 2032 1520 2112 1600
<< ptap >>
rect 0 0 2144 144
rect 0 1616 2144 1760
rect 0 0 144 1760
rect 2000 0 2144 1760
use LELOTR_RES4 XA1 
transform 1 0 280 0 1 280
box 280 280 1864 1480
<< labels >>
flabel metal1 s 16 16 2128 128 0 FreeSans 400 0 0 0 B
port 3 nsew signal bidirectional
flabel metal1 s 1534 1440 1930 1520 0 FreeSans 400 0 0 0 P
port 1 nsew signal bidirectional
flabel metal1 s 214 1440 610 1520 0 FreeSans 400 0 0 0 N
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2144 1760
<< end >>
