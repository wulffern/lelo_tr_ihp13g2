magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741993200
<< checkpaint >>
rect 0 0 152 152
<< metal1 >>
rect 0 0 152 152
<< via1 >>
rect 14 14 54 54
rect 14 98 54 138
rect 98 14 138 54
rect 98 98 138 138
<< metal2 >>
rect 0 0 152 152
<< via2 >>
rect 14 14 54 54
rect 14 98 54 138
rect 98 14 138 54
rect 98 98 138 138
<< metal3 >>
rect 0 0 152 152
<< via3 >>
rect 14 14 54 54
rect 14 98 54 138
rect 98 14 138 54
rect 98 98 138 138
<< metal4 >>
rect 0 0 152 152
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 152 152
<< end >>
