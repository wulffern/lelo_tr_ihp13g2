magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741993200
<< checkpaint >>
rect 0 0 1628 960
<< metal1 >>
rect 574 540 614 740
rect 1014 220 1054 420
rect 594 380 726 420
rect 726 860 1034 900
rect 726 380 766 900
rect 114 780 286 820
rect 114 260 546 300
rect 114 260 154 820
rect 506 220 594 260
rect 594 220 814 260
rect 814 540 1034 580
rect 814 220 854 580
rect 198 140 374 180
rect 198 460 374 500
rect 506 380 682 420
<< poly >>
rect 242 146 1386 174
rect 242 466 1386 494
rect 242 786 1386 814
<< metal4 >>
rect 946 0 1098 960
rect 506 0 658 960
rect 946 0 1098 960
rect 506 0 658 960
use LELOTR_NCHDL MN0 
transform 1 0 0 0 1 0
box 0 0 814 320
use LELOTR_NCHDL MN2 
transform 1 0 0 0 1 320
box 0 320 814 640
use LELOTR_NCHDL MN1 
transform 1 0 0 0 1 640
box 0 640 814 960
use LELOTR_PCHDL MP1 
transform 1 0 814 0 1 0
box 814 0 1628 320
use LELOTR_PCHDL MP0 
transform 1 0 814 0 1 320
box 814 320 1628 640
use LELOTR_PCHDL MP2 
transform 1 0 814 0 1 640
box 814 640 1628 960
use LELOTR_cut_M1M4_2x1 xcut0 
transform 1 0 946 0 1 60
box 946 60 1098 102
use LELOTR_cut_M1M4_2x1 xcut1 
transform 1 0 946 0 1 700
box 946 700 1098 742
use LELOTR_cut_M1M4_2x1 xcut2 
transform 1 0 506 0 1 60
box 506 60 658 102
use LELOTR_cut_M1M4_2x1 xcut3 
transform 1 0 506 0 1 860
box 506 860 658 902
<< labels >>
flabel metal1 s 198 140 374 180 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
flabel metal1 s 198 460 374 500 0 FreeSans 400 0 0 0 CK
port 2 nsew signal bidirectional
flabel metal1 s 506 380 682 420 0 FreeSans 400 0 0 0 Q
port 3 nsew signal bidirectional
flabel metal4 s 946 0 1098 960 0 FreeSans 400 0 0 0 AVDD
port 4 nsew signal bidirectional
flabel metal4 s 506 0 658 960 0 FreeSans 400 0 0 0 AVSS
port 5 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1628 960
<< end >>
